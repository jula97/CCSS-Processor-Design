module counter_6 (clk,clk2,clrn,clk3,out,segmentA,segmentB,segmentC,segmentD,segmentE,segmentF,segmentG); // a counter with 7-seg LED
input clk2,clrn; // clk, clear (active low)
input clk;
output clk3; // u==1: count up; u==0: count down
output [2:0] out; // 3-bit counter output
output segmentA, segmentB, segmentC, segmentD, segmentE, segmentF, segmentG; // seven-segment LED control
reg [2:0] out; // register type

clock_test_Clock_divider CLOCK(.clock_in(clk2), .clock_out(clk1));
assign clk3 = clk1;
always @ (posedge clk1 or negedge clrn) begin
//A Brief Introduction to Logic Circuits and Verilog HDL 59
if (!clrn) out <= 0; // if clrn is asserted, counter=0
else if (clk) out <= (out + 1) % 6; // if counter up, q++
//else if (q != 0) q <= q - 1; // else q–
//else out <= 4'd7;
end

bin27 display(
   .clk(clk1),
   .datain(out),
   .segmentA(segmentA),
   .segmentB(segmentB),
   .segmentC(segmentC),
   .segmentD(segmentD),
   .segmentE(segmentE),
   .segmentF(segmentF),
   .segmentG(segmentG) );
 
/* 
assign {g,f,e,d,c,b,a} = seg7(q); // call function to get LED control
function [6:0] seg7; // the function, 7-bit return value
input [2:0] q; // input argument
case (q) // cases:
3’d0 : seg7 = 7’b1000000; // 0’s LED control, 0: light on
3’d1 : seg7 = 7’b1111001; // 1’s LED control, 1: light off
3’d2 : seg7 = 7’b0100100; // 2’s LED control
3’d3 : seg7 = 7’b0110000; // 3’s LED control
3’d4 : seg7 = 7’b0011001; // 4’s LED control
3’d5 : seg7 = 7’b0010010; // 5’s LED control
default: seg7 = 7’b1111111; // default: all segments light off
endcase
endfunction*/

endmodule
